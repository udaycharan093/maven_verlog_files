review_uvm.sv
